library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
entity springdri is
port(con,en:in std_logic;
     spri:out std_logic_vector(0 to 1);
	  ligh:out std_logic_vector(0 to 2));
end entity springdri;
architecture behav of springdri is
begin
  beha:process(con,en)
  variable driver:std_logic_vector(0 to 4);
  variable cnt:std_logic_vector(7 downto 0);
  begin
    if en='0' then driver:="00000";
	 elsif con'event and con='1' then
	 cnt:=cnt+1;
		if    cnt="00000000" then driver:="01110";
		elsif cnt="00000001" then driver:="00100";
		elsif cnt="00000010" then driver:="11100";
		elsif cnt="00000011" then driver:="11111";
		elsif cnt="00000100" then driver:="10110";
		elsif cnt="00000101" then driver:="10000";
		elsif cnt="00000110" then driver:="10001";
		elsif cnt="00000111" then driver:="01011";
		elsif cnt="00001000" then driver:="11111";
		elsif cnt="00001001" then driver:="10001";
		elsif cnt="00001010" then driver:="01001";
		elsif cnt="00001011" then driver:="01010";
		elsif cnt="00001100" then driver:="00111";
		elsif cnt="00001101" then driver:="11001";
		elsif cnt="00001110" then driver:="10011";
		elsif cnt="00001111" then driver:="00011";
		elsif cnt="00010000" then driver:="10000";
		elsif cnt="00010001" then driver:="10001";
		elsif cnt="00010010" then driver:="11010";
		elsif cnt="00010011" then driver:="01011";
		elsif cnt="00010100" then driver:="10001";
		elsif cnt="00010101" then driver:="11101";
		elsif cnt="00010110" then driver:="01110";
		elsif cnt="00010111" then driver:="10111";
		elsif cnt="00011000" then driver:="00001";
		elsif cnt="00011001" then driver:="10111";
		elsif cnt="00011010" then driver:="11010";
		elsif cnt="00011011" then driver:="10000";
		elsif cnt="00011100" then driver:="01001";
		elsif cnt="00011101" then driver:="10011";
		elsif cnt="00011110" then driver:="11101";
		elsif cnt="00011111" then driver:="11010";
		elsif cnt="00100000" then driver:="01110";
		elsif cnt="00100001" then driver:="11111";
		elsif cnt="00100010" then driver:="00101";
		elsif cnt="00100011" then driver:="00011";
		elsif cnt="00100100" then driver:="01110";
		elsif cnt="00100101" then driver:="11110";
		elsif cnt="00100110" then driver:="10101";
		elsif cnt="00100111" then driver:="10011";
		elsif cnt="00101000" then driver:="11000";
		elsif cnt="00101001" then driver:="01101";
		elsif cnt="00101010" then driver:="11011";
		elsif cnt="00101011" then driver:="10101";
		elsif cnt="00101100" then driver:="10110";
		elsif cnt="00101101" then driver:="10101";
		elsif cnt="00101110" then driver:="10111";
		elsif cnt="00101111" then driver:="01101";
		elsif cnt="00110000" then driver:="01101";
		elsif cnt="00110001" then driver:="00001";
		elsif cnt="00110010" then driver:="11001";
		elsif cnt="00110011" then driver:="00001";
		elsif cnt="00110100" then driver:="00011";
		elsif cnt="00110101" then driver:="01001";
		elsif cnt="00110110" then driver:="01100";
		elsif cnt="00110111" then driver:="00111";
		elsif cnt="00111000" then driver:="10001";
		elsif cnt="00111001" then driver:="11010";
		elsif cnt="00111010" then driver:="10011";
		elsif cnt="00111011" then driver:="01100";
		elsif cnt="00111100" then driver:="10100";
		elsif cnt="00111101" then driver:="00001";
		elsif cnt="00111110" then driver:="10010";
		elsif cnt="00111111" then driver:="10101";
		elsif cnt="01000000" then driver:="11101";
		elsif cnt="01000001" then driver:="10101";
		elsif cnt="01000010" then driver:="01101";
		elsif cnt="01000011" then driver:="10100";
		elsif cnt="01000100" then driver:="01000";
		elsif cnt="01000101" then driver:="00010";
		elsif cnt="01000110" then driver:="01010";
		elsif cnt="01000111" then driver:="01110";
		elsif cnt="01001000" then driver:="11000";
		elsif cnt="01001001" then driver:="10101";
		elsif cnt="01001010" then driver:="10000";
		elsif cnt="01001011" then driver:="00001";
		elsif cnt="01001100" then driver:="11100";
		elsif cnt="01001101" then driver:="00010";
		elsif cnt="01001110" then driver:="11011";
		elsif cnt="01001111" then driver:="00101";
		elsif cnt="01010000" then driver:="10000";
		elsif cnt="01010001" then driver:="01111";
		elsif cnt="01010010" then driver:="11000";
		elsif cnt="01010011" then driver:="10110";
		elsif cnt="01010100" then driver:="00101";
		elsif cnt="01010101" then driver:="00110";
		elsif cnt="01010110" then driver:="11010";
		elsif cnt="01010111" then driver:="01001";
		elsif cnt="01011000" then driver:="00110";
		elsif cnt="01011001" then driver:="10000";
		elsif cnt="01011010" then driver:="01011";
		elsif cnt="01011011" then driver:="00100";
		elsif cnt="01011100" then driver:="00011";
		elsif cnt="01011101" then driver:="11001";
		elsif cnt="01011110" then driver:="01101";
		elsif cnt="01011111" then driver:="01110";
		elsif cnt="01100000" then driver:="10100";
		elsif cnt="01100001" then driver:="01011";
		elsif cnt="01100010" then driver:="00111";
		elsif cnt="01100011" then driver:="11100";
		elsif cnt="01100100" then driver:="00110";
		elsif cnt="01100101" then driver:="00110";
		elsif cnt="01100110" then driver:="00001";
		elsif cnt="01100111" then driver:="01011";
		elsif cnt="01101000" then driver:="01001";
		elsif cnt="01101001" then driver:="01000";
		elsif cnt="01101010" then driver:="10010";
		elsif cnt="01101011" then driver:="01101";
		elsif cnt="01101100" then driver:="00110";
		elsif cnt="01101101" then driver:="00011";
		elsif cnt="01101110" then driver:="10010";
		elsif cnt="01101111" then driver:="10011";
		elsif cnt="01110000" then driver:="10001";
		elsif cnt="01110001" then driver:="10001";
		elsif cnt="01110010" then driver:="11110";
		elsif cnt="01110011" then driver:="01010";
		elsif cnt="01110100" then driver:="00101";
		elsif cnt="01110101" then driver:="10100";
		elsif cnt="01110110" then driver:="10010";
		elsif cnt="01110111" then driver:="01110";
		elsif cnt="01111000" then driver:="00100";
		elsif cnt="01111001" then driver:="01111";
		elsif cnt="01111010" then driver:="10000";
		elsif cnt="01111011" then driver:="00110";
		elsif cnt="01111100" then driver:="11000";
		elsif cnt="01111101" then driver:="11101";
		elsif cnt="01111110" then driver:="00110";
		elsif cnt="01111111" then driver:="00101";
		elsif cnt="10000000" then driver:="10001";
		elsif cnt="10000001" then driver:="10001";
		elsif cnt="10000010" then driver:="00001";
		elsif cnt="10000011" then driver:="00011";
		elsif cnt="10000100" then driver:="01010";
		elsif cnt="10000101" then driver:="10001";
		elsif cnt="10000110" then driver:="11100";
		elsif cnt="10000111" then driver:="01100";
		elsif cnt="10001000" then driver:="11111";
		elsif cnt="10001001" then driver:="00110";
		elsif cnt="10001010" then driver:="01110";
		elsif cnt="10001011" then driver:="01100";
		elsif cnt="10001100" then driver:="11000";
		elsif cnt="10001101" then driver:="11001";
		elsif cnt="10001110" then driver:="01100";
		elsif cnt="10001111" then driver:="10010";
		elsif cnt="10010000" then driver:="11000";
		elsif cnt="10010001" then driver:="01000";
		elsif cnt="10010010" then driver:="11111";
		elsif cnt="10010011" then driver:="00100";
		elsif cnt="10010100" then driver:="10110";
		elsif cnt="10010101" then driver:="00101";
		elsif cnt="10010110" then driver:="11010";
		elsif cnt="10010111" then driver:="01001";
		elsif cnt="10011000" then driver:="00010";
		elsif cnt="10011001" then driver:="10011";
		elsif cnt="10011010" then driver:="01000";
		elsif cnt="10011011" then driver:="01110";
		elsif cnt="10011100" then driver:="01110";
		elsif cnt="10011101" then driver:="10111";
		elsif cnt="10011110" then driver:="10000";
		elsif cnt="10011111" then driver:="00100";
		elsif cnt="10100000" then driver:="11010";
		elsif cnt="10100001" then driver:="00100";
		elsif cnt="10100010" then driver:="01101";
		elsif cnt="10100011" then driver:="01110";
		elsif cnt="10100100" then driver:="01001";
		elsif cnt="10100101" then driver:="11110";
		elsif cnt="10100110" then driver:="01001";
		elsif cnt="10100111" then driver:="01101";
		elsif cnt="10101000" then driver:="01000";
		elsif cnt="10101001" then driver:="10111";
		elsif cnt="10101010" then driver:="00010";
		elsif cnt="10101011" then driver:="10101";
		elsif cnt="10101100" then driver:="01011";
		elsif cnt="10101101" then driver:="01101";
		elsif cnt="10101110" then driver:="11100";
		elsif cnt="10101111" then driver:="01100";
		elsif cnt="10110000" then driver:="10011";
		elsif cnt="10110001" then driver:="01111";
		elsif cnt="10110010" then driver:="00111";
		elsif cnt="10110011" then driver:="10100";
		elsif cnt="10110100" then driver:="11110";
		elsif cnt="10110101" then driver:="11011";
		elsif cnt="10110110" then driver:="00010";
		elsif cnt="10110111" then driver:="11010";
		elsif cnt="10111000" then driver:="01101";
		elsif cnt="10111001" then driver:="10110";
		elsif cnt="10111010" then driver:="11010";
		elsif cnt="10111011" then driver:="11000";
		elsif cnt="10111100" then driver:="10001";
		elsif cnt="10111101" then driver:="10011";
		elsif cnt="10111110" then driver:="01110";
		elsif cnt="10111111" then driver:="11111";
		elsif cnt="11000000" then driver:="01000";
		elsif cnt="11000001" then driver:="01100";
		elsif cnt="11000010" then driver:="10111";
		elsif cnt="11000011" then driver:="00010";
		elsif cnt="11000100" then driver:="11100";
		elsif cnt="11000101" then driver:="00011";
		elsif cnt="11000110" then driver:="01000";
		elsif cnt="11000111" then driver:="10000";
		elsif cnt="11001000" then driver:="01001";
		elsif cnt="11001001" then driver:="00010";
		elsif cnt="11001010" then driver:="00010";
		elsif cnt="11001011" then driver:="11111";
		elsif cnt="11001100" then driver:="00011";
		elsif cnt="11001101" then driver:="01101";
		elsif cnt="11001110" then driver:="01111";
		elsif cnt="11001111" then driver:="10001";
		elsif cnt="11010000" then driver:="01010";
		elsif cnt="11010001" then driver:="11111";
		elsif cnt="11010010" then driver:="11111";
		elsif cnt="11010011" then driver:="11101";
		elsif cnt="11010100" then driver:="10011";
		elsif cnt="11010101" then driver:="10001";
		elsif cnt="11010110" then driver:="00111";
		elsif cnt="11010111" then driver:="11111";
		elsif cnt="11011000" then driver:="00111";
		elsif cnt="11011001" then driver:="11101";
		elsif cnt="11011010" then driver:="01101";
		elsif cnt="11011011" then driver:="11011";
		elsif cnt="11011100" then driver:="00101";
		elsif cnt="11011101" then driver:="01111";
		elsif cnt="11011110" then driver:="01110";
		elsif cnt="11011111" then driver:="11011";
		elsif cnt="11100000" then driver:="10010";
		elsif cnt="11100001" then driver:="01110";
		elsif cnt="11100010" then driver:="10010";
		elsif cnt="11100011" then driver:="10001";
		elsif cnt="11100100" then driver:="10111";
		elsif cnt="11100101" then driver:="10001";
		elsif cnt="11100110" then driver:="11100";
		elsif cnt="11100111" then driver:="01110";
		elsif cnt="11101000" then driver:="11110";
		elsif cnt="11101001" then driver:="01110";
		elsif cnt="11101010" then driver:="11100";
		elsif cnt="11101011" then driver:="00101";
		elsif cnt="11101100" then driver:="10110";
		elsif cnt="11101101" then driver:="01010";
		elsif cnt="11101110" then driver:="11001";
		elsif cnt="11101111" then driver:="10100";
		elsif cnt="11110000" then driver:="01110";
		elsif cnt="11110001" then driver:="00010";
		elsif cnt="11110010" then driver:="00011";
		elsif cnt="11110011" then driver:="11100";
		elsif cnt="11110100" then driver:="10010";
		elsif cnt="11110101" then driver:="01101";
		elsif cnt="11110110" then driver:="11111";
		elsif cnt="11110111" then driver:="00010";
		elsif cnt="11111000" then driver:="10110";
		elsif cnt="11111001" then driver:="10000";
		elsif cnt="11111010" then driver:="00011";
		elsif cnt="11111011" then driver:="10111";
		elsif cnt="11111100" then driver:="01000";
		elsif cnt="11111101" then driver:="10110";
		elsif cnt="11111110" then driver:="10001";
		else                      driver:="11000";
		end if;
    end if;
	 spri <= driver(0 to 1);
	 ligh <= driver(2 to 4);
  end process beha;
end architecture behav;