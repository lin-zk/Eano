library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
entity vga_mode is
port(mode:in std_logic;
     clk0,clk1:in std_logic;
	  x0,y0,x1,y1: in integer range 0 to 200;
	  key:in std_logic_vector(0 to 20);
     vga_out_ram: in std_logic_vector(15 downto 0);
	  load:in std_logic;
     cho0,cho1:out std_logic;
	  vga_clk:buffer std_logic;
	  x,y:buffer integer range 0 to 200;
	  vga_out:out std_logic_vector(15 downto 0));
end entity vga_mode;
architecture behav of vga_mode is
signal chose:std_logic_vector(1 downto 0);
signal vga_out_tmp:std_logic_vector(15 downto 0);

constant key_w:std_logic_vector(15 downto 0):=x"FFFF";
constant key_b:std_logic_vector(15 downto 0):=x"0000";
constant key_c:std_logic_vector(15 downto 0):=x"E7FF";
begin
  chose <= "10" when mode='1'else
           "01" when mode='0'else
			  "00";
  cho0 <= chose(0);
  cho1 <= chose(1);
  vga_clk <= clk1 when mode='1'else
             clk0 when mode='0'else
			    '0';
  y <= y1+3 when mode='1'else
       y0 when mode='0'else
		 0;
  x <= x1 when mode='1'else
       x0 when mode='0'else
		 0;
rdcl:process(x,y)
  begin
    if load='1'then
	   if y<=90 then
		  if y>=30 and y<=57 then
		    if x>=35 and x<=123 then
				if x=35 and y=33 then vga_out_tmp <= x"0000";
				elsif x=36 and y=33 then vga_out_tmp <= x"0000";
				elsif x=37 and y=33 then vga_out_tmp <= x"0000";
				elsif x=38 and y=33 then vga_out_tmp <= x"0000";
				elsif x=39 and y=33 then vga_out_tmp <= x"0000";
				elsif x=40 and y=33 then vga_out_tmp <= x"0000";
				elsif x=41 and y=33 then vga_out_tmp <= x"0000";
				elsif x=42 and y=33 then vga_out_tmp <= x"0000";
				elsif x=43 and y=33 then vga_out_tmp <= x"0000";
				elsif x=44 and y=33 then vga_out_tmp <= x"0000";
				elsif x=45 and y=33 then vga_out_tmp <= x"0000";
				elsif x=46 and y=33 then vga_out_tmp <= x"0000";
				elsif x=47 and y=33 then vga_out_tmp <= x"0000";
				elsif x=48 and y=33 then vga_out_tmp <= x"0000";
				elsif x=37 and y=34 then vga_out_tmp <= x"0000";
				elsif x=38 and y=34 then vga_out_tmp <= x"0000";
				elsif x=39 and y=34 then vga_out_tmp <= x"0000";
				elsif x=40 and y=34 then vga_out_tmp <= x"0000";
				elsif x=44 and y=34 then vga_out_tmp <= x"0000";
				elsif x=45 and y=34 then vga_out_tmp <= x"0000";
				elsif x=46 and y=34 then vga_out_tmp <= x"0000";
				elsif x=47 and y=34 then vga_out_tmp <= x"0000";
				elsif x=48 and y=34 then vga_out_tmp <= x"0000";
				elsif x=49 and y=34 then vga_out_tmp <= x"0000";
				elsif x=37 and y=35 then vga_out_tmp <= x"0000";
				elsif x=38 and y=35 then vga_out_tmp <= x"0000";
				elsif x=39 and y=35 then vga_out_tmp <= x"0000";
				elsif x=40 and y=35 then vga_out_tmp <= x"0000";
				elsif x=46 and y=35 then vga_out_tmp <= x"0000";
				elsif x=47 and y=35 then vga_out_tmp <= x"0000";
				elsif x=48 and y=35 then vga_out_tmp <= x"0000";
				elsif x=49 and y=35 then vga_out_tmp <= x"0000";
				elsif x=37 and y=36 then vga_out_tmp <= x"0000";
				elsif x=38 and y=36 then vga_out_tmp <= x"0000";
				elsif x=39 and y=36 then vga_out_tmp <= x"0000";
				elsif x=40 and y=36 then vga_out_tmp <= x"0000";
				elsif x=47 and y=36 then vga_out_tmp <= x"0000";
				elsif x=48 and y=36 then vga_out_tmp <= x"0000";
				elsif x=49 and y=36 then vga_out_tmp <= x"0000";
				elsif x=37 and y=37 then vga_out_tmp <= x"0000";
				elsif x=38 and y=37 then vga_out_tmp <= x"0000";
				elsif x=39 and y=37 then vga_out_tmp <= x"0000";
				elsif x=40 and y=37 then vga_out_tmp <= x"0000";
				elsif x=48 and y=37 then vga_out_tmp <= x"0000";
				elsif x=49 and y=37 then vga_out_tmp <= x"0000";
				elsif x=37 and y=38 then vga_out_tmp <= x"0000";
				elsif x=38 and y=38 then vga_out_tmp <= x"0000";
				elsif x=39 and y=38 then vga_out_tmp <= x"0000";
				elsif x=40 and y=38 then vga_out_tmp <= x"0000";
				elsif x=37 and y=39 then vga_out_tmp <= x"0000";
				elsif x=38 and y=39 then vga_out_tmp <= x"0000";
				elsif x=39 and y=39 then vga_out_tmp <= x"0000";
				elsif x=40 and y=39 then vga_out_tmp <= x"0000";
				elsif x=45 and y=39 then vga_out_tmp <= x"0000";
				elsif x=46 and y=39 then vga_out_tmp <= x"0000";
				elsif x=37 and y=40 then vga_out_tmp <= x"0000";
				elsif x=38 and y=40 then vga_out_tmp <= x"0000";
				elsif x=39 and y=40 then vga_out_tmp <= x"0000";
				elsif x=40 and y=40 then vga_out_tmp <= x"0000";
				elsif x=45 and y=40 then vga_out_tmp <= x"0000";
				elsif x=46 and y=40 then vga_out_tmp <= x"0000";
				elsif x=62 and y=40 then vga_out_tmp <= x"0000";
				elsif x=63 and y=40 then vga_out_tmp <= x"0000";
				elsif x=64 and y=40 then vga_out_tmp <= x"0000";
				elsif x=65 and y=40 then vga_out_tmp <= x"0000";
				elsif x=66 and y=40 then vga_out_tmp <= x"0000";
				elsif x=67 and y=40 then vga_out_tmp <= x"0000";
				elsif x=68 and y=40 then vga_out_tmp <= x"0000";
				elsif x=69 and y=40 then vga_out_tmp <= x"0000";
				elsif x=70 and y=40 then vga_out_tmp <= x"0000";
				elsif x=83 and y=40 then vga_out_tmp <= x"0000";
				elsif x=84 and y=40 then vga_out_tmp <= x"0000";
				elsif x=85 and y=40 then vga_out_tmp <= x"0000";
				elsif x=86 and y=40 then vga_out_tmp <= x"0000";
				elsif x=87 and y=40 then vga_out_tmp <= x"0000";
				elsif x=89 and y=40 then vga_out_tmp <= x"0000";
				elsif x=90 and y=40 then vga_out_tmp <= x"0000";
				elsif x=91 and y=40 then vga_out_tmp <= x"0000";
				elsif x=92 and y=40 then vga_out_tmp <= x"0000";
				elsif x=93 and y=40 then vga_out_tmp <= x"0000";
				elsif x=94 and y=40 then vga_out_tmp <= x"0000";
				elsif x=95 and y=40 then vga_out_tmp <= x"0000";
				elsif x=111 and y=40 then vga_out_tmp <= x"0000";
				elsif x=112 and y=40 then vga_out_tmp <= x"0000";
				elsif x=113 and y=40 then vga_out_tmp <= x"0000";
				elsif x=114 and y=40 then vga_out_tmp <= x"0000";
				elsif x=115 and y=40 then vga_out_tmp <= x"0000";
				elsif x=116 and y=40 then vga_out_tmp <= x"0000";
				elsif x=117 and y=40 then vga_out_tmp <= x"0000";
				elsif x=118 and y=40 then vga_out_tmp <= x"0000";
				elsif x=37 and y=41 then vga_out_tmp <= x"0000";
				elsif x=38 and y=41 then vga_out_tmp <= x"0000";
				elsif x=39 and y=41 then vga_out_tmp <= x"0000";
				elsif x=40 and y=41 then vga_out_tmp <= x"0000";
				elsif x=45 and y=41 then vga_out_tmp <= x"0000";
				elsif x=46 and y=41 then vga_out_tmp <= x"0000";
				elsif x=61 and y=41 then vga_out_tmp <= x"0000";
				elsif x=62 and y=41 then vga_out_tmp <= x"0000";
				elsif x=63 and y=41 then vga_out_tmp <= x"0000";
				elsif x=64 and y=41 then vga_out_tmp <= x"0000";
				elsif x=65 and y=41 then vga_out_tmp <= x"0000";
				elsif x=67 and y=41 then vga_out_tmp <= x"0000";
				elsif x=68 and y=41 then vga_out_tmp <= x"0000";
				elsif x=69 and y=41 then vga_out_tmp <= x"0000";
				elsif x=70 and y=41 then vga_out_tmp <= x"0000";
				elsif x=71 and y=41 then vga_out_tmp <= x"0000";
				elsif x=83 and y=41 then vga_out_tmp <= x"0000";
				elsif x=84 and y=41 then vga_out_tmp <= x"0000";
				elsif x=85 and y=41 then vga_out_tmp <= x"0000";
				elsif x=86 and y=41 then vga_out_tmp <= x"0000";
				elsif x=87 and y=41 then vga_out_tmp <= x"0000";
				elsif x=88 and y=41 then vga_out_tmp <= x"0000";
				elsif x=89 and y=41 then vga_out_tmp <= x"0000";
				elsif x=90 and y=41 then vga_out_tmp <= x"0000";
				elsif x=91 and y=41 then vga_out_tmp <= x"0000";
				elsif x=92 and y=41 then vga_out_tmp <= x"0000";
				elsif x=93 and y=41 then vga_out_tmp <= x"0000";
				elsif x=94 and y=41 then vga_out_tmp <= x"0000";
				elsif x=95 and y=41 then vga_out_tmp <= x"0000";
				elsif x=110 and y=41 then vga_out_tmp <= x"0000";
				elsif x=111 and y=41 then vga_out_tmp <= x"0000";
				elsif x=112 and y=41 then vga_out_tmp <= x"0000";
				elsif x=113 and y=41 then vga_out_tmp <= x"0000";
				elsif x=114 and y=41 then vga_out_tmp <= x"0000";
				elsif x=115 and y=41 then vga_out_tmp <= x"0000";
				elsif x=116 and y=41 then vga_out_tmp <= x"0000";
				elsif x=117 and y=41 then vga_out_tmp <= x"0000";
				elsif x=118 and y=41 then vga_out_tmp <= x"0000";
				elsif x=119 and y=41 then vga_out_tmp <= x"0000";
				elsif x=37 and y=42 then vga_out_tmp <= x"0000";
				elsif x=38 and y=42 then vga_out_tmp <= x"0000";
				elsif x=39 and y=42 then vga_out_tmp <= x"0000";
				elsif x=40 and y=42 then vga_out_tmp <= x"0000";
				elsif x=44 and y=42 then vga_out_tmp <= x"0000";
				elsif x=45 and y=42 then vga_out_tmp <= x"0000";
				elsif x=46 and y=42 then vga_out_tmp <= x"0000";
				elsif x=60 and y=42 then vga_out_tmp <= x"0000";
				elsif x=61 and y=42 then vga_out_tmp <= x"0000";
				elsif x=62 and y=42 then vga_out_tmp <= x"0000";
				elsif x=63 and y=42 then vga_out_tmp <= x"0000";
				elsif x=69 and y=42 then vga_out_tmp <= x"0000";
				elsif x=70 and y=42 then vga_out_tmp <= x"0000";
				elsif x=71 and y=42 then vga_out_tmp <= x"0000";
				elsif x=85 and y=42 then vga_out_tmp <= x"0000";
				elsif x=86 and y=42 then vga_out_tmp <= x"0000";
				elsif x=87 and y=42 then vga_out_tmp <= x"0000";
				elsif x=88 and y=42 then vga_out_tmp <= x"0000";
				elsif x=89 and y=42 then vga_out_tmp <= x"0000";
				elsif x=93 and y=42 then vga_out_tmp <= x"0000";
				elsif x=94 and y=42 then vga_out_tmp <= x"0000";
				elsif x=95 and y=42 then vga_out_tmp <= x"0000";
				elsif x=96 and y=42 then vga_out_tmp <= x"0000";
				elsif x=109 and y=42 then vga_out_tmp <= x"0000";
				elsif x=110 and y=42 then vga_out_tmp <= x"0000";
				elsif x=111 and y=42 then vga_out_tmp <= x"0000";
				elsif x=112 and y=42 then vga_out_tmp <= x"0000";
				elsif x=117 and y=42 then vga_out_tmp <= x"0000";
				elsif x=118 and y=42 then vga_out_tmp <= x"0000";
				elsif x=119 and y=42 then vga_out_tmp <= x"0000";
				elsif x=120 and y=42 then vga_out_tmp <= x"0000";
				elsif x=37 and y=43 then vga_out_tmp <= x"0000";
				elsif x=38 and y=43 then vga_out_tmp <= x"0000";
				elsif x=39 and y=43 then vga_out_tmp <= x"0000";
				elsif x=40 and y=43 then vga_out_tmp <= x"0000";
				elsif x=41 and y=43 then vga_out_tmp <= x"0000";
				elsif x=42 and y=43 then vga_out_tmp <= x"0000";
				elsif x=43 and y=43 then vga_out_tmp <= x"0000";
				elsif x=44 and y=43 then vga_out_tmp <= x"0000";
				elsif x=45 and y=43 then vga_out_tmp <= x"0000";
				elsif x=46 and y=43 then vga_out_tmp <= x"0000";
				elsif x=60 and y=43 then vga_out_tmp <= x"0000";
				elsif x=61 and y=43 then vga_out_tmp <= x"0000";
				elsif x=62 and y=43 then vga_out_tmp <= x"0000";
				elsif x=63 and y=43 then vga_out_tmp <= x"0000";
				elsif x=69 and y=43 then vga_out_tmp <= x"0000";
				elsif x=70 and y=43 then vga_out_tmp <= x"0000";
				elsif x=71 and y=43 then vga_out_tmp <= x"0000";
				elsif x=72 and y=43 then vga_out_tmp <= x"0000";
				elsif x=85 and y=43 then vga_out_tmp <= x"0000";
				elsif x=86 and y=43 then vga_out_tmp <= x"0000";
				elsif x=87 and y=43 then vga_out_tmp <= x"0000";
				elsif x=88 and y=43 then vga_out_tmp <= x"0000";
				elsif x=94 and y=43 then vga_out_tmp <= x"0000";
				elsif x=95 and y=43 then vga_out_tmp <= x"0000";
				elsif x=96 and y=43 then vga_out_tmp <= x"0000";
				elsif x=109 and y=43 then vga_out_tmp <= x"0000";
				elsif x=110 and y=43 then vga_out_tmp <= x"0000";
				elsif x=111 and y=43 then vga_out_tmp <= x"0000";
				elsif x=118 and y=43 then vga_out_tmp <= x"0000";
				elsif x=119 and y=43 then vga_out_tmp <= x"0000";
				elsif x=120 and y=43 then vga_out_tmp <= x"0000";
				elsif x=37 and y=44 then vga_out_tmp <= x"0000";
				elsif x=38 and y=44 then vga_out_tmp <= x"0000";
				elsif x=39 and y=44 then vga_out_tmp <= x"0000";
				elsif x=40 and y=44 then vga_out_tmp <= x"0000";
				elsif x=43 and y=44 then vga_out_tmp <= x"0000";
				elsif x=44 and y=44 then vga_out_tmp <= x"0000";
				elsif x=45 and y=44 then vga_out_tmp <= x"0000";
				elsif x=46 and y=44 then vga_out_tmp <= x"0000";
				elsif x=61 and y=44 then vga_out_tmp <= x"0000";
				elsif x=62 and y=44 then vga_out_tmp <= x"0000";
				elsif x=63 and y=44 then vga_out_tmp <= x"0000";
				elsif x=69 and y=44 then vga_out_tmp <= x"0000";
				elsif x=70 and y=44 then vga_out_tmp <= x"0000";
				elsif x=71 and y=44 then vga_out_tmp <= x"0000";
				elsif x=72 and y=44 then vga_out_tmp <= x"0000";
				elsif x=85 and y=44 then vga_out_tmp <= x"0000";
				elsif x=86 and y=44 then vga_out_tmp <= x"0000";
				elsif x=87 and y=44 then vga_out_tmp <= x"0000";
				elsif x=94 and y=44 then vga_out_tmp <= x"0000";
				elsif x=95 and y=44 then vga_out_tmp <= x"0000";
				elsif x=96 and y=44 then vga_out_tmp <= x"0000";
				elsif x=108 and y=44 then vga_out_tmp <= x"0000";
				elsif x=109 and y=44 then vga_out_tmp <= x"0000";
				elsif x=110 and y=44 then vga_out_tmp <= x"0000";
				elsif x=111 and y=44 then vga_out_tmp <= x"0000";
				elsif x=118 and y=44 then vga_out_tmp <= x"0000";
				elsif x=119 and y=44 then vga_out_tmp <= x"0000";
				elsif x=120 and y=44 then vga_out_tmp <= x"0000";
				elsif x=121 and y=44 then vga_out_tmp <= x"0000";
				elsif x=37 and y=45 then vga_out_tmp <= x"0000";
				elsif x=38 and y=45 then vga_out_tmp <= x"0000";
				elsif x=39 and y=45 then vga_out_tmp <= x"0000";
				elsif x=40 and y=45 then vga_out_tmp <= x"0000";
				elsif x=45 and y=45 then vga_out_tmp <= x"0000";
				elsif x=46 and y=45 then vga_out_tmp <= x"0000";
				elsif x=66 and y=45 then vga_out_tmp <= x"0000";
				elsif x=67 and y=45 then vga_out_tmp <= x"0000";
				elsif x=68 and y=45 then vga_out_tmp <= x"0000";
				elsif x=69 and y=45 then vga_out_tmp <= x"0000";
				elsif x=70 and y=45 then vga_out_tmp <= x"0000";
				elsif x=71 and y=45 then vga_out_tmp <= x"0000";
				elsif x=72 and y=45 then vga_out_tmp <= x"0000";
				elsif x=85 and y=45 then vga_out_tmp <= x"0000";
				elsif x=86 and y=45 then vga_out_tmp <= x"0000";
				elsif x=87 and y=45 then vga_out_tmp <= x"0000";
				elsif x=94 and y=45 then vga_out_tmp <= x"0000";
				elsif x=95 and y=45 then vga_out_tmp <= x"0000";
				elsif x=96 and y=45 then vga_out_tmp <= x"0000";
				elsif x=108 and y=45 then vga_out_tmp <= x"0000";
				elsif x=109 and y=45 then vga_out_tmp <= x"0000";
				elsif x=110 and y=45 then vga_out_tmp <= x"0000";
				elsif x=111 and y=45 then vga_out_tmp <= x"0000";
				elsif x=119 and y=45 then vga_out_tmp <= x"0000";
				elsif x=120 and y=45 then vga_out_tmp <= x"0000";
				elsif x=121 and y=45 then vga_out_tmp <= x"0000";
				elsif x=37 and y=46 then vga_out_tmp <= x"0000";
				elsif x=38 and y=46 then vga_out_tmp <= x"0000";
				elsif x=39 and y=46 then vga_out_tmp <= x"0000";
				elsif x=40 and y=46 then vga_out_tmp <= x"0000";
				elsif x=45 and y=46 then vga_out_tmp <= x"0000";
				elsif x=46 and y=46 then vga_out_tmp <= x"0000";
				elsif x=63 and y=46 then vga_out_tmp <= x"0000";
				elsif x=64 and y=46 then vga_out_tmp <= x"0000";
				elsif x=65 and y=46 then vga_out_tmp <= x"0000";
				elsif x=66 and y=46 then vga_out_tmp <= x"0000";
				elsif x=67 and y=46 then vga_out_tmp <= x"0000";
				elsif x=68 and y=46 then vga_out_tmp <= x"0000";
				elsif x=69 and y=46 then vga_out_tmp <= x"0000";
				elsif x=70 and y=46 then vga_out_tmp <= x"0000";
				elsif x=71 and y=46 then vga_out_tmp <= x"0000";
				elsif x=72 and y=46 then vga_out_tmp <= x"0000";
				elsif x=85 and y=46 then vga_out_tmp <= x"0000";
				elsif x=86 and y=46 then vga_out_tmp <= x"0000";
				elsif x=87 and y=46 then vga_out_tmp <= x"0000";
				elsif x=94 and y=46 then vga_out_tmp <= x"0000";
				elsif x=95 and y=46 then vga_out_tmp <= x"0000";
				elsif x=96 and y=46 then vga_out_tmp <= x"0000";
				elsif x=108 and y=46 then vga_out_tmp <= x"0000";
				elsif x=109 and y=46 then vga_out_tmp <= x"0000";
				elsif x=110 and y=46 then vga_out_tmp <= x"0000";
				elsif x=119 and y=46 then vga_out_tmp <= x"0000";
				elsif x=120 and y=46 then vga_out_tmp <= x"0000";
				elsif x=121 and y=46 then vga_out_tmp <= x"0000";
				elsif x=37 and y=47 then vga_out_tmp <= x"0000";
				elsif x=38 and y=47 then vga_out_tmp <= x"0000";
				elsif x=39 and y=47 then vga_out_tmp <= x"0000";
				elsif x=40 and y=47 then vga_out_tmp <= x"0000";
				elsif x=45 and y=47 then vga_out_tmp <= x"0000";
				elsif x=46 and y=47 then vga_out_tmp <= x"0000";
				elsif x=61 and y=47 then vga_out_tmp <= x"0000";
				elsif x=62 and y=47 then vga_out_tmp <= x"0000";
				elsif x=63 and y=47 then vga_out_tmp <= x"0000";
				elsif x=64 and y=47 then vga_out_tmp <= x"0000";
				elsif x=65 and y=47 then vga_out_tmp <= x"0000";
				elsif x=66 and y=47 then vga_out_tmp <= x"0000";
				elsif x=69 and y=47 then vga_out_tmp <= x"0000";
				elsif x=70 and y=47 then vga_out_tmp <= x"0000";
				elsif x=71 and y=47 then vga_out_tmp <= x"0000";
				elsif x=72 and y=47 then vga_out_tmp <= x"0000";
				elsif x=85 and y=47 then vga_out_tmp <= x"0000";
				elsif x=86 and y=47 then vga_out_tmp <= x"0000";
				elsif x=87 and y=47 then vga_out_tmp <= x"0000";
				elsif x=94 and y=47 then vga_out_tmp <= x"0000";
				elsif x=95 and y=47 then vga_out_tmp <= x"0000";
				elsif x=96 and y=47 then vga_out_tmp <= x"0000";
				elsif x=108 and y=47 then vga_out_tmp <= x"0000";
				elsif x=109 and y=47 then vga_out_tmp <= x"0000";
				elsif x=110 and y=47 then vga_out_tmp <= x"0000";
				elsif x=119 and y=47 then vga_out_tmp <= x"0000";
				elsif x=120 and y=47 then vga_out_tmp <= x"0000";
				elsif x=121 and y=47 then vga_out_tmp <= x"0000";
				elsif x=37 and y=48 then vga_out_tmp <= x"0000";
				elsif x=38 and y=48 then vga_out_tmp <= x"0000";
				elsif x=39 and y=48 then vga_out_tmp <= x"0000";
				elsif x=40 and y=48 then vga_out_tmp <= x"0000";
				elsif x=60 and y=48 then vga_out_tmp <= x"0000";
				elsif x=61 and y=48 then vga_out_tmp <= x"0000";
				elsif x=62 and y=48 then vga_out_tmp <= x"0000";
				elsif x=63 and y=48 then vga_out_tmp <= x"0000";
				elsif x=64 and y=48 then vga_out_tmp <= x"0000";
				elsif x=69 and y=48 then vga_out_tmp <= x"0000";
				elsif x=70 and y=48 then vga_out_tmp <= x"0000";
				elsif x=71 and y=48 then vga_out_tmp <= x"0000";
				elsif x=72 and y=48 then vga_out_tmp <= x"0000";
				elsif x=85 and y=48 then vga_out_tmp <= x"0000";
				elsif x=86 and y=48 then vga_out_tmp <= x"0000";
				elsif x=87 and y=48 then vga_out_tmp <= x"0000";
				elsif x=94 and y=48 then vga_out_tmp <= x"0000";
				elsif x=95 and y=48 then vga_out_tmp <= x"0000";
				elsif x=96 and y=48 then vga_out_tmp <= x"0000";
				elsif x=108 and y=48 then vga_out_tmp <= x"0000";
				elsif x=109 and y=48 then vga_out_tmp <= x"0000";
				elsif x=110 and y=48 then vga_out_tmp <= x"0000";
				elsif x=119 and y=48 then vga_out_tmp <= x"0000";
				elsif x=120 and y=48 then vga_out_tmp <= x"0000";
				elsif x=121 and y=48 then vga_out_tmp <= x"0000";
				elsif x=37 and y=49 then vga_out_tmp <= x"0000";
				elsif x=38 and y=49 then vga_out_tmp <= x"0000";
				elsif x=39 and y=49 then vga_out_tmp <= x"0000";
				elsif x=40 and y=49 then vga_out_tmp <= x"0000";
				elsif x=49 and y=49 then vga_out_tmp <= x"0000";
				elsif x=50 and y=49 then vga_out_tmp <= x"0000";
				elsif x=60 and y=49 then vga_out_tmp <= x"0000";
				elsif x=61 and y=49 then vga_out_tmp <= x"0000";
				elsif x=62 and y=49 then vga_out_tmp <= x"0000";
				elsif x=63 and y=49 then vga_out_tmp <= x"0000";
				elsif x=69 and y=49 then vga_out_tmp <= x"0000";
				elsif x=70 and y=49 then vga_out_tmp <= x"0000";
				elsif x=71 and y=49 then vga_out_tmp <= x"0000";
				elsif x=72 and y=49 then vga_out_tmp <= x"0000";
				elsif x=85 and y=49 then vga_out_tmp <= x"0000";
				elsif x=86 and y=49 then vga_out_tmp <= x"0000";
				elsif x=87 and y=49 then vga_out_tmp <= x"0000";
				elsif x=94 and y=49 then vga_out_tmp <= x"0000";
				elsif x=95 and y=49 then vga_out_tmp <= x"0000";
				elsif x=96 and y=49 then vga_out_tmp <= x"0000";
				elsif x=108 and y=49 then vga_out_tmp <= x"0000";
				elsif x=109 and y=49 then vga_out_tmp <= x"0000";
				elsif x=110 and y=49 then vga_out_tmp <= x"0000";
				elsif x=119 and y=49 then vga_out_tmp <= x"0000";
				elsif x=120 and y=49 then vga_out_tmp <= x"0000";
				elsif x=121 and y=49 then vga_out_tmp <= x"0000";
				elsif x=37 and y=50 then vga_out_tmp <= x"0000";
				elsif x=38 and y=50 then vga_out_tmp <= x"0000";
				elsif x=39 and y=50 then vga_out_tmp <= x"0000";
				elsif x=40 and y=50 then vga_out_tmp <= x"0000";
				elsif x=48 and y=50 then vga_out_tmp <= x"0000";
				elsif x=49 and y=50 then vga_out_tmp <= x"0000";
				elsif x=50 and y=50 then vga_out_tmp <= x"0000";
				elsif x=60 and y=50 then vga_out_tmp <= x"0000";
				elsif x=61 and y=50 then vga_out_tmp <= x"0000";
				elsif x=62 and y=50 then vga_out_tmp <= x"0000";
				elsif x=69 and y=50 then vga_out_tmp <= x"0000";
				elsif x=70 and y=50 then vga_out_tmp <= x"0000";
				elsif x=71 and y=50 then vga_out_tmp <= x"0000";
				elsif x=72 and y=50 then vga_out_tmp <= x"0000";
				elsif x=85 and y=50 then vga_out_tmp <= x"0000";
				elsif x=86 and y=50 then vga_out_tmp <= x"0000";
				elsif x=87 and y=50 then vga_out_tmp <= x"0000";
				elsif x=94 and y=50 then vga_out_tmp <= x"0000";
				elsif x=95 and y=50 then vga_out_tmp <= x"0000";
				elsif x=96 and y=50 then vga_out_tmp <= x"0000";
				elsif x=108 and y=50 then vga_out_tmp <= x"0000";
				elsif x=109 and y=50 then vga_out_tmp <= x"0000";
				elsif x=110 and y=50 then vga_out_tmp <= x"0000";
				elsif x=111 and y=50 then vga_out_tmp <= x"0000";
				elsif x=118 and y=50 then vga_out_tmp <= x"0000";
				elsif x=119 and y=50 then vga_out_tmp <= x"0000";
				elsif x=120 and y=50 then vga_out_tmp <= x"0000";
				elsif x=121 and y=50 then vga_out_tmp <= x"0000";
				elsif x=37 and y=51 then vga_out_tmp <= x"0000";
				elsif x=38 and y=51 then vga_out_tmp <= x"0000";
				elsif x=39 and y=51 then vga_out_tmp <= x"0000";
				elsif x=40 and y=51 then vga_out_tmp <= x"0000";
				elsif x=48 and y=51 then vga_out_tmp <= x"0000";
				elsif x=49 and y=51 then vga_out_tmp <= x"0000";
				elsif x=60 and y=51 then vga_out_tmp <= x"0000";
				elsif x=61 and y=51 then vga_out_tmp <= x"0000";
				elsif x=62 and y=51 then vga_out_tmp <= x"0000";
				elsif x=69 and y=51 then vga_out_tmp <= x"0000";
				elsif x=70 and y=51 then vga_out_tmp <= x"0000";
				elsif x=71 and y=51 then vga_out_tmp <= x"0000";
				elsif x=72 and y=51 then vga_out_tmp <= x"0000";
				elsif x=73 and y=51 then vga_out_tmp <= x"0000";
				elsif x=74 and y=51 then vga_out_tmp <= x"0000";
				elsif x=85 and y=51 then vga_out_tmp <= x"0000";
				elsif x=86 and y=51 then vga_out_tmp <= x"0000";
				elsif x=87 and y=51 then vga_out_tmp <= x"0000";
				elsif x=94 and y=51 then vga_out_tmp <= x"0000";
				elsif x=95 and y=51 then vga_out_tmp <= x"0000";
				elsif x=96 and y=51 then vga_out_tmp <= x"0000";
				elsif x=108 and y=51 then vga_out_tmp <= x"0000";
				elsif x=109 and y=51 then vga_out_tmp <= x"0000";
				elsif x=110 and y=51 then vga_out_tmp <= x"0000";
				elsif x=111 and y=51 then vga_out_tmp <= x"0000";
				elsif x=118 and y=51 then vga_out_tmp <= x"0000";
				elsif x=119 and y=51 then vga_out_tmp <= x"0000";
				elsif x=120 and y=51 then vga_out_tmp <= x"0000";
				elsif x=121 and y=51 then vga_out_tmp <= x"0000";
				elsif x=37 and y=52 then vga_out_tmp <= x"0000";
				elsif x=38 and y=52 then vga_out_tmp <= x"0000";
				elsif x=39 and y=52 then vga_out_tmp <= x"0000";
				elsif x=40 and y=52 then vga_out_tmp <= x"0000";
				elsif x=47 and y=52 then vga_out_tmp <= x"0000";
				elsif x=48 and y=52 then vga_out_tmp <= x"0000";
				elsif x=49 and y=52 then vga_out_tmp <= x"0000";
				elsif x=60 and y=52 then vga_out_tmp <= x"0000";
				elsif x=61 and y=52 then vga_out_tmp <= x"0000";
				elsif x=62 and y=52 then vga_out_tmp <= x"0000";
				elsif x=63 and y=52 then vga_out_tmp <= x"0000";
				elsif x=68 and y=52 then vga_out_tmp <= x"0000";
				elsif x=69 and y=52 then vga_out_tmp <= x"0000";
				elsif x=70 and y=52 then vga_out_tmp <= x"0000";
				elsif x=71 and y=52 then vga_out_tmp <= x"0000";
				elsif x=72 and y=52 then vga_out_tmp <= x"0000";
				elsif x=73 and y=52 then vga_out_tmp <= x"0000";
				elsif x=74 and y=52 then vga_out_tmp <= x"0000";
				elsif x=85 and y=52 then vga_out_tmp <= x"0000";
				elsif x=86 and y=52 then vga_out_tmp <= x"0000";
				elsif x=87 and y=52 then vga_out_tmp <= x"0000";
				elsif x=94 and y=52 then vga_out_tmp <= x"0000";
				elsif x=95 and y=52 then vga_out_tmp <= x"0000";
				elsif x=96 and y=52 then vga_out_tmp <= x"0000";
				elsif x=109 and y=52 then vga_out_tmp <= x"0000";
				elsif x=110 and y=52 then vga_out_tmp <= x"0000";
				elsif x=111 and y=52 then vga_out_tmp <= x"0000";
				elsif x=112 and y=52 then vga_out_tmp <= x"0000";
				elsif x=117 and y=52 then vga_out_tmp <= x"0000";
				elsif x=118 and y=52 then vga_out_tmp <= x"0000";
				elsif x=119 and y=52 then vga_out_tmp <= x"0000";
				elsif x=120 and y=52 then vga_out_tmp <= x"0000";
				elsif x=37 and y=53 then vga_out_tmp <= x"0000";
				elsif x=38 and y=53 then vga_out_tmp <= x"0000";
				elsif x=39 and y=53 then vga_out_tmp <= x"0000";
				elsif x=40 and y=53 then vga_out_tmp <= x"0000";
				elsif x=44 and y=53 then vga_out_tmp <= x"0000";
				elsif x=45 and y=53 then vga_out_tmp <= x"0000";
				elsif x=46 and y=53 then vga_out_tmp <= x"0000";
				elsif x=47 and y=53 then vga_out_tmp <= x"0000";
				elsif x=48 and y=53 then vga_out_tmp <= x"0000";
				elsif x=49 and y=53 then vga_out_tmp <= x"0000";
				elsif x=60 and y=53 then vga_out_tmp <= x"0000";
				elsif x=61 and y=53 then vga_out_tmp <= x"0000";
				elsif x=62 and y=53 then vga_out_tmp <= x"0000";
				elsif x=63 and y=53 then vga_out_tmp <= x"0000";
				elsif x=64 and y=53 then vga_out_tmp <= x"0000";
				elsif x=66 and y=53 then vga_out_tmp <= x"0000";
				elsif x=67 and y=53 then vga_out_tmp <= x"0000";
				elsif x=68 and y=53 then vga_out_tmp <= x"0000";
				elsif x=69 and y=53 then vga_out_tmp <= x"0000";
				elsif x=70 and y=53 then vga_out_tmp <= x"0000";
				elsif x=71 and y=53 then vga_out_tmp <= x"0000";
				elsif x=72 and y=53 then vga_out_tmp <= x"0000";
				elsif x=73 and y=53 then vga_out_tmp <= x"0000";
				elsif x=74 and y=53 then vga_out_tmp <= x"0000";
				elsif x=85 and y=53 then vga_out_tmp <= x"0000";
				elsif x=86 and y=53 then vga_out_tmp <= x"0000";
				elsif x=87 and y=53 then vga_out_tmp <= x"0000";
				elsif x=88 and y=53 then vga_out_tmp <= x"0000";
				elsif x=93 and y=53 then vga_out_tmp <= x"0000";
				elsif x=94 and y=53 then vga_out_tmp <= x"0000";
				elsif x=95 and y=53 then vga_out_tmp <= x"0000";
				elsif x=96 and y=53 then vga_out_tmp <= x"0000";
				elsif x=97 and y=53 then vga_out_tmp <= x"0000";
				elsif x=110 and y=53 then vga_out_tmp <= x"0000";
				elsif x=111 and y=53 then vga_out_tmp <= x"0000";
				elsif x=112 and y=53 then vga_out_tmp <= x"0000";
				elsif x=113 and y=53 then vga_out_tmp <= x"0000";
				elsif x=114 and y=53 then vga_out_tmp <= x"0000";
				elsif x=115 and y=53 then vga_out_tmp <= x"0000";
				elsif x=116 and y=53 then vga_out_tmp <= x"0000";
				elsif x=117 and y=53 then vga_out_tmp <= x"0000";
				elsif x=118 and y=53 then vga_out_tmp <= x"0000";
				elsif x=119 and y=53 then vga_out_tmp <= x"0000";
				elsif x=35 and y=54 then vga_out_tmp <= x"0000";
				elsif x=36 and y=54 then vga_out_tmp <= x"0000";
				elsif x=37 and y=54 then vga_out_tmp <= x"0000";
				elsif x=38 and y=54 then vga_out_tmp <= x"0000";
				elsif x=39 and y=54 then vga_out_tmp <= x"0000";
				elsif x=40 and y=54 then vga_out_tmp <= x"0000";
				elsif x=41 and y=54 then vga_out_tmp <= x"0000";
				elsif x=42 and y=54 then vga_out_tmp <= x"0000";
				elsif x=43 and y=54 then vga_out_tmp <= x"0000";
				elsif x=44 and y=54 then vga_out_tmp <= x"0000";
				elsif x=45 and y=54 then vga_out_tmp <= x"0000";
				elsif x=46 and y=54 then vga_out_tmp <= x"0000";
				elsif x=47 and y=54 then vga_out_tmp <= x"0000";
				elsif x=48 and y=54 then vga_out_tmp <= x"0000";
				elsif x=49 and y=54 then vga_out_tmp <= x"0000";
				elsif x=61 and y=54 then vga_out_tmp <= x"0000";
				elsif x=62 and y=54 then vga_out_tmp <= x"0000";
				elsif x=63 and y=54 then vga_out_tmp <= x"0000";
				elsif x=64 and y=54 then vga_out_tmp <= x"0000";
				elsif x=65 and y=54 then vga_out_tmp <= x"0000";
				elsif x=66 and y=54 then vga_out_tmp <= x"0000";
				elsif x=67 and y=54 then vga_out_tmp <= x"0000";
				elsif x=68 and y=54 then vga_out_tmp <= x"0000";
				elsif x=70 and y=54 then vga_out_tmp <= x"0000";
				elsif x=71 and y=54 then vga_out_tmp <= x"0000";
				elsif x=72 and y=54 then vga_out_tmp <= x"0000";
				elsif x=73 and y=54 then vga_out_tmp <= x"0000";
				elsif x=74 and y=54 then vga_out_tmp <= x"0000";
				elsif x=83 and y=54 then vga_out_tmp <= x"0000";
				elsif x=84 and y=54 then vga_out_tmp <= x"0000";
				elsif x=85 and y=54 then vga_out_tmp <= x"0000";
				elsif x=86 and y=54 then vga_out_tmp <= x"0000";
				elsif x=87 and y=54 then vga_out_tmp <= x"0000";
				elsif x=88 and y=54 then vga_out_tmp <= x"0000";
				elsif x=89 and y=54 then vga_out_tmp <= x"0000";
				elsif x=92 and y=54 then vga_out_tmp <= x"0000";
				elsif x=93 and y=54 then vga_out_tmp <= x"0000";
				elsif x=94 and y=54 then vga_out_tmp <= x"0000";
				elsif x=95 and y=54 then vga_out_tmp <= x"0000";
				elsif x=96 and y=54 then vga_out_tmp <= x"0000";
				elsif x=97 and y=54 then vga_out_tmp <= x"0000";
				elsif x=98 and y=54 then vga_out_tmp <= x"0000";
				elsif x=111 and y=54 then vga_out_tmp <= x"0000";
				elsif x=112 and y=54 then vga_out_tmp <= x"0000";
				elsif x=113 and y=54 then vga_out_tmp <= x"0000";
				elsif x=114 and y=54 then vga_out_tmp <= x"0000";
				elsif x=115 and y=54 then vga_out_tmp <= x"0000";
				elsif x=116 and y=54 then vga_out_tmp <= x"0000";
				elsif x=117 and y=54 then vga_out_tmp <= x"0000";
				elsif x=118 and y=54 then vga_out_tmp <= x"0000";
				else vga_out_tmp<=x"FFFF";
				end if;
			 end if;
	     elsif x<20 then
		    vga_out_tmp <= x"FFFF";
		  elsif x<2*20 then
		    vga_out_tmp <= x"F800";
		  elsif x<3*20 then
		    vga_out_tmp <= x"F5E3";
		  elsif x<4*20 then
		    vga_out_tmp <= x"FFE0";
		  elsif x<5*20 then
		    vga_out_tmp <= x"07EF";
		  elsif x<6*20 then
		    vga_out_tmp <= x"07FF";
		  elsif x<7*20 then
		    vga_out_tmp <= x"867D";
		  elsif x<8*20 then
		    vga_out_tmp <= x"8010";
		  else
		    vga_out_tmp <= x"481F";
		  end if;
		else
		  vga_out_tmp <= x"0000";
		end if;
	 else
      if y>25 then
        if x>= 7 and x<=153 then
		    if x<=7*2-1 then 
		      if key(0)='1' then vga_out_tmp <= key_c;
			   else vga_out_tmp <= key_w;
			   end if;
		    elsif x <= 7*3-1 then 
		      if key(1)='1' then vga_out_tmp <= key_c;
			   else vga_out_tmp <= key_b;
			   end if;
		    elsif x <= 7*4-1 then 
		      if key(2)='1' then vga_out_tmp <= key_c;
			   else vga_out_tmp <= key_w;
			   end if;
		    elsif x <= 7*5-1 then
		      if key(3)='1' then vga_out_tmp <= key_c;
			   else vga_out_tmp <= key_b;
			   end if;
		    elsif x <= 7*6-1 then
		      if key(4)='1' then vga_out_tmp <= key_c;
			   else vga_out_tmp <= key_w;
			   end if;
		    elsif x <= 7*7-1 then
		      if key(5)='1' then vga_out_tmp <= key_c;
			   else vga_out_tmp <= key_b;
			   end if;
		    elsif x <= 7*8-1 then
		      if key(6)='1' then vga_out_tmp <= key_c;
			   else vga_out_tmp <= key_w;
			   end if;
		    elsif x <= 7*9-1 then
		      if key(7)='1' then vga_out_tmp <= key_c;
			   else vga_out_tmp <= key_b;
			   end if;
		    elsif x <= 7*10-1 then
		      if key(8)='1' then vga_out_tmp <= key_c;
			   else vga_out_tmp <= key_w;
			   end if;
		    elsif x <= 7*11-1 then
		      if key(9)='1' then vga_out_tmp <= key_c;
			   else vga_out_tmp <= key_b;
			   end if;
		    elsif x <= 7*12-1 then
		      if key(10)='1' then vga_out_tmp <= key_c;
			   else vga_out_tmp <= key_w;
			   end if;
		    elsif x <= 7*13-1 then
		      if key(11)='1' then vga_out_tmp <= key_c;
			   else vga_out_tmp <= key_b;
			   end if;
		    elsif x <= 7*14-1 then
		      if key(12)='1' then vga_out_tmp <= key_c;
			   else vga_out_tmp <= key_w;
			   end if;
		    elsif x <= 7*15-1 then
		      if key(13)='1' then vga_out_tmp <= key_c;
			   else vga_out_tmp <= key_b;
			   end if;
		    elsif x <= 7*16-1 then
		      if key(14)='1' then vga_out_tmp <= key_c;
			   else vga_out_tmp <= key_w;
			   end if;
		    elsif x <= 7*17-1 then
		      if key(15)='1' then vga_out_tmp <= key_c;
			   else vga_out_tmp <= key_b;
			   end if;
		    elsif x <= 7*18-1 then
		      if key(16)='1' then vga_out_tmp <= key_c;
			   else vga_out_tmp <= key_w;
			   end if;
		    elsif x <= 7*19-1 then
		      if key(17)='1' then vga_out_tmp <= key_c;
			   else vga_out_tmp <= key_b;
			   end if;
		    elsif x <= 7*20-1 then
		      if key(18)='1' then vga_out_tmp <= key_c;
			   else vga_out_tmp <= key_w;
			   end if;
		    elsif x <= 7*21-1 then
		      if key(19)='1' then vga_out_tmp <= key_c;
			   else vga_out_tmp <= key_b;
			   end if;
		    else
		      if key(20)='1' then vga_out_tmp <= key_c;
			   else vga_out_tmp <= key_w;
			   end if;
		    end if;
		  else vga_out_tmp <= vga_out_ram;
	     end if;
	    else vga_out_tmp <= vga_out_ram;
      end if;
	 end if;
  end process rdcl;
vout:process(vga_clk)
  begin
    if vga_clk'event and vga_clk='1' then
      vga_out <= vga_out_tmp;
    end if;
  end process vout;
end architecture behav;
