library ieee;
use ieee.std_logic_1164.all;
entity SEG_datactrl is
port(space,enter,esc,load:in std_logic;
     music:in std_logic_vector(0 to 20);
     d0,d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17:
	  out std_logic_vector(5 downto 0));
end entity SEG_datactrl;
architecture behav of SEG_datactrl is
begin
  process(space,enter,esc,load,music)
    begin
	 if load='1' then --Loading...
	   d0 <= "010101";
		d1 <= "011000";
		d2 <= "001010";
		d3 <= "001101";
		d4 <= "010010";
		d5 <= "010111";
		d6 <= "010000";
		d7 <= "111110";
		d8 <= "111110";
		d9 <= "111110";
		d10 <= "000000";
		d11 <= "000000";
		d12 <= "000000";
		d13 <= "111111";
	 elsif esc='1' then--SATING...
	   d0 <= "011100";
		d1 <= "001010";
		d2 <= "011101";
		d3 <= "010010";
		d4 <= "010111";
		d5 <= "010000";
		d6 <= "111110";
		d7 <= "111110";
		d8 <= "111110";
		d9 <= "000000";
		d10 <= "000000";
		d11 <= "000000";
		d12 <= "111111";
		d13 <= "111111";
	 elsif enter='1' then--RESET
	   d0 <= "011011";
		d1 <= "001110";
		d2 <= "011100";
		d3 <= "011101";
		d4 <= "001010";
		d5 <= "111111";
		d6 <= "111111";
		d7 <= "111111";
		d8 <= "111111";
		d9 <= "111111";
		d10 <= "111111";
		d11 <= "111111";
		d12 <= "111111";
		d13 <= "111111";
	 elsif space='1' then--STOPING...
	   d0 <= "011100";
		d1 <= "011101";
		d2 <= "011000";
		d3 <= "011001";
		d4 <= "010010";
		d5 <= "010111";
		d6 <= "010000";
		d7 <= "000000";
		d8 <= "000000";
		d9 <= "000000";
		d10 <= "111111";
		d11 <= "111111";
		d12 <= "111111";
		d13 <= "111111";
	 elsif music/="000000000000000000000" then--PLAYING...
	   d0 <= "011001";
		d1 <= "010101";
		d2 <= "001010";
		d3 <= "100010";
		d4 <= "010010";
		d5 <= "010111";
		d6 <= "010000";
		d7 <= "111110";
		d8 <= "111110";
		d9 <= "111110";
		d10 <= "000000"; 
		d11 <= "000000";
		d12 <= "000000";
		d13 <= "111111";
	 else --HEllo.EANO
	   d0 <= "010001";
	   d1 <= "101000";
      d2 <= "000001";
      d3 <= "000001";
      d4 <= "110010";
      d5 <= "111110";
      d6 <= "001110";
      d7 <= "001010";
      d8 <= "010111";
      d9 <= "011000";
      d10 <= "000000";
      d11 <= "000000";
      d12 <= "000000";
      d13 <= "111111";
	 end if;
  end process;
end architecture behav;